--
-- cgrom.vhd
--
-- MZ-700 CG-ROM pattern module
-- for MZ-700 on FPGA
--
-- Nibbles Lab. 2005
--

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

--  Uncomment the following lines to use the declarations that are
--  provided for instantiating Xilinx primitive components.
library UNISIM;
use UNISIM.VComponents.all;

entity cgrom is
    Port ( ROMA : in std_logic_vector(10 downto 0);
           CSEL : in std_logic;
           ROMD : out std_logic_vector(7 downto 0);
		 PCGSW : in std_logic;
		 CSPCG : in std_logic;
		 WR : in std_logic;
           RAMA : in std_logic_vector(1 downto 0);
           RAMD : in std_logic_vector(7 downto 0);
		 MCLK : in std_logic;
		 DCLK : in std_logic);
end cgrom;

architecture Behavioral of cgrom is

--
-- CG-ROM
--
signal net_gnd : std_logic_vector(7 downto 0);
signal net_vcc : std_logic;
signal XA : std_logic_vector(10 downto 0);
signal D0 : std_logic_vector(7 downto 0);
signal D1 : std_logic_vector(7 downto 0);
signal CPYD0 : std_logic_vector(7 downto 0);
signal CPYD1 : std_logic_vector(7 downto 0);
--
-- PCG
--
signal EXA : std_logic_vector(10 downto 0);
signal D2 : std_logic_vector(7 downto 0);
signal CPYA : std_logic_vector(10 downto 0);
signal PCGA : std_logic_vector(10 downto 0);
signal TMPA : std_logic_vector(2 downto 0);
signal BUFD : std_logic_vector(7 downto 0);
signal PCGD : std_logic_vector(7 downto 0);
signal PCGWP : std_logic;
signal PCGDSEL : std_logic;
signal TMPDSEL : std_logic;

begin

	--
	-- fixed signals
	--
	net_gnd<=(others=>'0');
	net_vcc<='1';
	--
	-- reverse address signal
	--
	XA<=ROMA(10 downto 5)&(not ROMA(4 downto 0));
	EXA<=CSEL&XA(9 downto 0);

	--
	-- Font select
	--
	process( CSEL, XA(10), PCGSW, D0, D1, D2 ) begin
		if( CSEL='0' ) then
			if( PCGSW='0' ) then
				ROMD<=D0;
			else
				if( XA(10)='0' ) then
					ROMD<=D0;
				else
					ROMD<=D2;
				end if;
			end if;
		else
			if( PCGSW='0' ) then
				ROMD<=D1;
			else
				if( XA(10)='0' ) then
					ROMD<=D1;
				else
					ROMD<=D2;
				end if;
			end if;
		end if;
	end process;

	--
	-- Access Registers
	--
	process( MCLK ) begin
		if( MCLK'event and MCLK='1' ) then
			PCGA(10 downto 8)<=TMPA;
			PCGDSEL<=TMPDSEL;
			if( CSPCG='0' and WR='0' ) then
				if( RAMA="00" ) then
					BUFD<=RAMD;
				elsif( RAMA="01" ) then
					PCGA(7 downto 0)<=RAMD(7 downto 5)&(not RAMD(4 downto 0));
				elsif( RAMA="10" ) then
					TMPA<=RAMD(2 downto 0);
					PCGWP<=not RAMD(4);
					TMPDSEL<=RAMD(5);
				end if;
			end if;
		end if;
	end process;
	CPYA<='1'&TMPA(1 downto 0)&PCGA(7 downto 0);
	PCGD<=BUFD when PCGDSEL='0' else
		 CPYD0 when PCGDSEL='1' and PCGA(10)='0' else
		 CPYD1;

	--
	-- RAM (CG data included:normal)
	--
   RAMB16_S9_S9_inst0 : RAMB16_S9_S9
	generic map (
      INIT_A => X"000", --  Value of output RAM registers on Port A at startup
      INIT_B => X"000", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"000", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"000", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "READ_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "READ_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
		INIT_00 => X"00000000000000001824427E424242007C22223C22227C001C22404040221C00",
		INIT_01 => X"78242222222478007E40407840407E007E404078404040001C22404E42221C00",
		INIT_02 => X"4242427E424242001C08080808081C000E040404044438004244487048444200",
		INIT_03 => X"4040404040407E0042665A5A424242004262524A464242001824424242241800",
		INIT_04 => X"7C42427C40404000182442424A241A007C42427C484442003C42403C02423C00",
		INIT_05 => X"3E080808080808004242424242423C0042424224241818004242425A5A664200",
		INIT_06 => X"42422418244242002222221C080808007E02041820407E0008080808FF080808",
		INIT_07 => X"080808080F00000008080808F8000000080808080F08080808080808FF000000",
		INIT_08 => X"3C42465A62423C000818280808083E003C42020C30407E003C42023C02423C00",
		INIT_09 => X"040C14247E0404007E407804024438001C20407C42423C007E42040810101000",
		INIT_0A => X"3C42423C42423C003C42423E020438000000007E0000000000007E007E000000",
		INIT_0B => X"0000080000080810000204081020400000000000001818000000000000080810",
		INIT_0C => X"00FF000000000000404040404040404080808080808080FF01010101010101FF",
		INIT_0D => X"000000FF000000001010101010101010FFFF000000000000C0C0C0C0C0C0C0C0",
		INIT_0E => X"0000000000FF0000040404040404040400000000FFFFFFFF0F0F0F0F0F0F0F0F",
		INIT_0F => X"00000000000000FF0101010101010101000000000000FFFF0303030303030303",
		INIT_10 => X"00000804FE040800081C3E7F7F1C3E00FF7F3F1F0F070301FFFFFFFFFFFFFFFF",
		INIT_11 => X"081C3E7F3E1C0800000010207F201000081C2A7F2A080800003C7E7E7E7E3C00",
		INIT_12 => X"003C424242423C003C42020C10001000FFC381818181C3FF0000000003040808",
		INIT_13 => X"00000000C020101080C0E0F0F8FCFEFF0103070F1F3F7FFF0000080000080000",
		INIT_14 => X"00081C2A080808000E18306030180E003C20202020203C00367F7F7F3E1C0800",
		INIT_15 => X"3C04040404043C001C224A564C201E00FFFEFCF8F0E0C08070180C060C187000",
		INIT_16 => X"A050A050A050A0500040201008040200AA55AA55AA55AA55F0F0F0F00F0F0F0F",
		INIT_17 => X"000000000F08080800000000F808080808080808F808080800000000FF080808",
		INIT_18 => X"0000013E541414000808080800000800242424000000000024247E247E242400",
		INIT_19 => X"081E281C0A3C08000062640810264600304848304A443A000408100000000000",
		INIT_1A => X"040810101008040020100808081020000008083E08080000082A1C3E1C2A0800",
		INIT_1B => X"0F0F0F0FF0F0F0F08142241818244281101020C0000000000808040300000000",
		INIT_1C => X"FF000000000000008080808080808080FF80808080808080FF01010101010101",
		INIT_1D => X"0000FF0000000000202020202020202001020408102040808040201008040201",
		INIT_1E => X"00000000FF0000000808080808080808FFFFFFFF00000000F0F0F0F0F0F0F0F0",
		INIT_1F => X"000000000000FF0002020202020202020000000000FFFFFF0707070707070707",
		INIT_20 => X"000808082A1C08000438083E08081000003E020202023E000022221202041800",
		INIT_21 => X"003002320204380002040818280808000008042222222200083E083E08080800",
		INIT_22 => X"001E122202041800001C000000003E00003E0202140804000404040404081000",
		INIT_23 => X"2424242404081000003E103E10100E00001C001C003C02001C003E0202040800",
		INIT_24 => X"103E121410100E00001E122A06041800003E0204081422001010101814101000",
		INIT_25 => X"103E12121212240008083E080810200020203E2020201E001C003E0808081000",
		INIT_26 => X"143E1414040810000030000202043800002A2A2A02040800003E222222223E00",
		INIT_27 => X"101E2404040408001E1010100000000000003E020C0810000000103E12141000",
		INIT_28 => X"003E222202040800003E021408142000003E0202020418003E020A0C08081000",
		INIT_29 => X"083E222202040800003E080808083E00043E040C1424040010103E1214101000",
		INIT_2A => X"001C040404043E00003E023E02023E00083E08082A2A08000010280402020000",
		INIT_2B => X"00202022242830000002021408142000000828282A2A2C00083E04081C2A0800",
		INIT_2C => X"00081020223E0200000000080808780000000408182808000000001C04043E00",
		INIT_2D => X"003E023E0204080000000000402010000000083E22020C0000003C043C043C00",
		INIT_2E => X"705070000000000000000000000020000000003E08083E000000002A2A020C00",
		INIT_2F => X"104820000000000000000000705070000000043E0C1424000000001C00000000",
		INIT_30 => X"1C1C3E1C08003E00FFF7F7F7D5E3F7FFFFF7E3D5F7F7F7FFFFFFF7FB81FBF7FF",
		INIT_31 => X"FFFFEFDF81DFEFFFBBBBBB83BBBBBBFFE3DDBFBFBFDDE3FF18247EFF5A240000",
		INIT_32 => X"E047427E4247E000223E2A0808497F411C1C083E080814220011D2FCD2110000",
		INIT_33 => X"00884B3F4B880000221408083E081C1C3C7EFFDBFFE77E3C3C4281A58199423C",
		INIT_34 => X"3E22223E22223E003E223E223E224200082A2A081422410008093A0C1C2A4900",
		INIT_35 => X"08083E081C2A490008143E493E1C7F000008083E08087F0008487E483E087F00",
		INIT_36 => X"203E483C287E0800047E547F527F0A000814227F1212240038127F173B521400",
		INIT_37 => X"7F49497F4141410022143E083E0808000C12103810103E0000C0C85454552200",
		INIT_38 => X"000000000002FF020202020202020702020202020202FF020000205088050200",
		INIT_39 => X"000E1122C404020100FF008142428100007088442320408000C4A4948F94A4C4",
		INIT_3A => X"00232529F12925238890A0C0C0A898B8A8B0B8C0C0A09088804020101F204080",
		INIT_3B => X"00002424E724240008083E00003E0808081020100804020455AA55AA55AA55AA",
		INIT_3C => X"0000000000000000007070700000000000070707000000000077777700000000",
		INIT_3D => X"0000000000707070007070700070707000070707007070700077777700707070",
		INIT_3E => X"0000000000070707007070700007070700070707000707070077777700070707",
		INIT_3F => X"0000000000777777007070700077777700070707007777770077777700777777",
		INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
	port map (
      DOA => D0,      -- Port A 8-bit Data Output
      DOB => CPYD0,      -- Port B 8-bit Data Output
      DOPA => open,    -- Port A 1-bit Parity Output
      DOPB => open,    -- Port B 1-bit Parity Output
      ADDRA => XA,  -- Port A 11-bit Address Input
      ADDRB => CPYA,  -- Port B 11-bit Address Input
      CLKA => DCLK,    -- Port A Clock
      CLKB => PCGDSEL,    -- Port B Clock
      DIA => net_gnd,      -- Port A 8-bit Data Input
      DIB => net_gnd,      -- Port B 8-bit Data Input
      DIPA => net_gnd(0 downto 0),    -- Port A 1-bit parity Input
      DIPB => net_gnd(0 downto 0),    -- Port-B 1-bit parity Input
      ENA => net_vcc,      -- Port A RAM Enable Input
      ENB => net_vcc,      -- PortB RAM Enable Input
      SSRA => net_gnd(0),    -- Port A Synchronous Set/Reset Input
      SSRB => net_gnd(0),    -- Port B Synchronous Set/Reset Input
      WEA => net_gnd(0),      -- Port A Write Enable Input
      WEB => net_gnd(0)       -- Port B Write Enable Input
	);

	--
	-- RAM (CG data included:alternate)
	--
   RAMB16_S9_S9_inst1 : RAMB16_S9_S9
	generic map (
      INIT_A => X"000", --  Value of output RAM registers on Port A at startup
      INIT_B => X"000", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"000", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"000", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "READ_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "READ_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
		INIT_00 => X"0000000000000000000038043C443A0040405C6242625C0000003C4240423C00",
		INIT_01 => X"02023A4642463A0000003C427E403C000C12107C1010100000003A46463A023C",
		INIT_02 => X"40405C62424242000800180808081C0004000C04040444384040444850684400",
		INIT_03 => X"1808080808081C00000076494949490000005C624242420000003C4242423C00",
		INIT_04 => X"00005C62625C404000003A46463A020200005C624040400000003E403C027C00",
		INIT_05 => X"10107C1010120C000000424242423C0000004242422418000000414949493600",
		INIT_06 => X"000044281028440000004242463A023C00007E0418207E0008080808FF080808",
		INIT_07 => X"080808080F00000008080808F8000000080808080F08080808080808FF000000",
		INIT_08 => X"3C42465A62423C000818280808083E003C42020C30407E003C42023C02423C00",
		INIT_09 => X"040C14247E0404007E407804024438001C20407C42423C007E42040810101000",
		INIT_0A => X"3C42423C42423C003C42423E020438000000007E0000000000007E007E000000",
		INIT_0B => X"0000080000080810000204081020400000000000001818000000000000080810",
		INIT_0C => X"00FF000000000000404040404040404080808080808080FF01010101010101FF",
		INIT_0D => X"000000FF000000001010101010101010FFFF000000000000C0C0C0C0C0C0C0C0",
		INIT_0E => X"0000000000FF0000040404040404040400000000FFFFFFFF0F0F0F0F0F0F0F0F",
		INIT_0F => X"00000000000000FF0101010101010101000000000000FFFF0303030303030303",
		INIT_10 => X"00000804FE040800081C3E7F7F1C3E00FF7F3F1F0F070301FFFFFFFFFFFFFFFF",
		INIT_11 => X"081C3E7F3E1C0800000010207F201000081C2A7F2A080800003C7E7E7E7E3C00",
		INIT_12 => X"003C424242423C003C42020C10001000FFC381818181C3FF0000000003040808",
		INIT_13 => X"00000000C020101080C0E0F0F8FCFEFF0103070F1F3F7FFF0000080000080000",
		INIT_14 => X"00081C2A080808000E18306030180E003C20202020203C00367F7F7F3E1C0800",
		INIT_15 => X"3C04040404043C001C224A564C201E00FFFEFCF8F0E0C08070180C060C187000",
		INIT_16 => X"A050A050A050A0500040201008040200AA55AA55AA55AA55F0F0F0F00F0F0F0F",
		INIT_17 => X"000000000F08080800000000F808080808080808F808080800000000FF080808",
		INIT_18 => X"0000013E541414000808080800000800242424000000000024247E247E242400",
		INIT_19 => X"081E281C0A3C08000062640810264600304848304A443A000408100000000000",
		INIT_1A => X"040810101008040020100808081020000008083E08080000082A1C3E1C2A0800",
		INIT_1B => X"0F0F0F0FF0F0F0F08142241818244281101020C0000000000808040300000000",
		INIT_1C => X"FF000000000000008080808080808080FF80808080808080FF01010101010101",
		INIT_1D => X"0000FF0000000000202020202020202004081122448810202010884422110804",
		INIT_1E => X"00000000FF0000000808080808080808FFFFFFFF00000000F0F0F0F0F0F0F0F0",
		INIT_1F => X"000000000000FF0002020202020202020000000000FFFFFF0707070707070707",
		INIT_20 => X"000808082A1C080010FE207C0202FC0000FC020000807E003C08107E08100C00",
		INIT_21 => X"40404040444438008482828282906000849E84849CA65C00107E087E04026018",
		INIT_22 => X"0C18306030180C009E8080808090DE00107E107E10709C723854929292926400",
		INIT_23 => X"444444640408100020F820F822221C007010147E9494640060009CA2C2821C00",
		INIT_24 => X"4444FE4458403E0020FC405E80A0BE0008FE08384838081020222C3040807E00",
		INIT_25 => X"22F925242424480020FA41449CA61C00E026458484887000FE04081010080400",
		INIT_26 => X"20FE1008442018001020207048888600807C0202020418007C08102C42022418",
		INIT_27 => X"84BE8484848448001E101010000000000020702078946800000058E428201000",
		INIT_28 => X"20E42A3262A2240004447C4AB29766003800104A4A8A300020FC207CAA926400",
		INIT_29 => X"18003C420204080010007C081028460020FD217CA2A26400484C32E224101008",
		INIT_2A => X"089CAACACA8C1800080E0808788E78009E849E849CA6DC000020508804020200",
		INIT_2B => X"20E62C3464A4220004447C4AB29264007C08103C421A241820E42A3266AB2600",
		INIT_2C => X"20FD2160A0623E0000000000080808780000484444442000000010B8D4983000",
		INIT_2D => X"10FE2074B8487E00000000000040201000200078040408000000203820786000",
		INIT_2E => X"705070000000000000000000000020000020007810304C00000000F804041800",
		INIT_2F => X"209040000000000000000000007050700020742078A468000000001C00000000",
		INIT_30 => X"1C1C3E1C08003E00FFF7F7F7D5E3F7FFFFF7E3D5F7F7F7FFFFFFF7FB81FBF7FF",
		INIT_31 => X"FFFFEFDF81DFEFFFBBBBBB83BBBBBBFFE3DDBFBFBFDDE3FF18247EFF5A240000",
		INIT_32 => X"E047427E4247E000223E2A0808497F411C1C083E080814220011D2FCD2110000",
		INIT_33 => X"00884B3F4B880000221408083E081C1C3C7EFFDBFFE77E3C3C4281A58199423C",
		INIT_34 => X"3E22223E22223E003E223E223E224200082A2A081422410008093A0C1C2A4900",
		INIT_35 => X"08083E081C2A490008143E493E1C7F000008083E08087F0008487E483E087F00",
		INIT_36 => X"203E483C287E0800047E547F527F0A000814227F1212240038127F173B521400",
		INIT_37 => X"7F49497F4141410022143E083E0808000C12103810103E0000C0C85454552200",
		INIT_38 => X"000000000002FF020202020202020702020202020202FF020000205088050200",
		INIT_39 => X"000E1122C404020100FF008142428100007088442320408000C4A4948F94A4C4",
		INIT_3A => X"00232529F12925238890A0C0C0A898B8A8B0B8C0C0A09088804020101F204080",
		INIT_3B => X"00002424E724240008083E00003E0808081020100804020455AA55AA55AA55AA",
		INIT_3C => X"0000000000000000007070700000000000070707000000000077777700000000",
		INIT_3D => X"0000000000707070007070700070707000070707007070700077777700707070",
		INIT_3E => X"0000000000070707007070700007070700070707000707070077777700070707",
		INIT_3F => X"0000000000777777007070700077777700070707007777770077777700777777",
		INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
	port map (
      DOA => D1,      -- Port A 8-bit Data Output
      DOB => CPYD1,      -- Port B 8-bit Data Output
      DOPA => open,    -- Port A 1-bit Parity Output
      DOPB => open,    -- Port B 1-bit Parity Output
      ADDRA => XA,  -- Port A 11-bit Address Input
      ADDRB => CPYA,  -- Port B 11-bit Address Input
      CLKA => DCLK,    -- Port A Clock
      CLKB => PCGDSEL,    -- Port B Clock
      DIA => net_gnd,      -- Port A 8-bit Data Input
      DIB => net_gnd,      -- Port B 8-bit Data Input
      DIPA => net_gnd(0 downto 0),    -- Port A 1-bit parity Input
      DIPB => net_gnd(0 downto 0),    -- Port-B 1-bit parity Input
      ENA => net_vcc,      -- Port A RAM Enable Input
      ENB => net_vcc,      -- PortB RAM Enable Input
      SSRA => net_gnd(0),    -- Port A Synchronous Set/Reset Input
      SSRB => net_gnd(0),    -- Port B Synchronous Set/Reset Input
      WEA => net_gnd(0),      -- Port A Write Enable Input
      WEB => net_gnd(0)       -- Port B Write Enable Input
	);

	--
	-- RAM (PCG data area)
	--
   RAMB16_S9_S9_inst2 : RAMB16_S9_S9
   generic map (
      INIT_A => X"000", --  Value of output RAM registers on Port A at startup
      INIT_B => X"000", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"000", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"000", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "READ_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "READ_FIRST") --  WRITE_FIRST, READ_FIRST or NO_CHANGE
   port map (
      DOA => D2,      -- Port A 8-bit Data Output
      DOB => open,      -- Port B 8-bit Data Output
      DOPA => open,    -- Port A 1-bit Parity Output
      DOPB => open,    -- Port B 1-bit Parity Output
      ADDRA => EXA,  -- Port A 11-bit Address Input
      ADDRB => PCGA,  -- Port B 11-bit Address Input
      CLKA => DCLK,    -- Port A Clock
      CLKB => PCGWP,    -- Port B Clock
      DIA => net_gnd,      -- Port A 8-bit Data Input
      DIB => PCGD,      -- Port B 8-bit Data Input
      DIPA => net_gnd(0 downto 0),    -- Port A 1-bit parity Input
      DIPB => net_gnd(0 downto 0),    -- Port-B 1-bit parity Input
      ENA => net_vcc,      -- Port A RAM Enable Input
      ENB => net_vcc,      -- PortB RAM Enable Input
      SSRA => net_gnd(0),    -- Port A Synchronous Set/Reset Input
      SSRB => net_gnd(0),    -- Port B Synchronous Set/Reset Input
      WEA => net_gnd(0),      -- Port A Write Enable Input
      WEB => net_vcc       -- Port B Write Enable Input
   );

end Behavioral;
