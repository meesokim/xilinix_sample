--
-- mom.vhd
--
-- MONITOR 1Z-009A/MZ NEW-MONITOR module
-- for MZ-700 on FPGA
--
-- Nibbles Lab. 2005
--

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

--  Uncomment the following lines to use the declarations that are
--  provided for instantiating Xilinx primitive components.
library UNISIM;
use UNISIM.VComponents.all;

entity mrom is
    Port ( A : in std_logic_vector(11 downto 0);
           CS : in std_logic;
           D : out std_logic_vector(7 downto 0);
		 CLK : in std_logic);
end mrom;

architecture Behavioral of mrom is

--
-- signals
--
signal net_gnd : std_logic_vector(7 downto 0);
signal net_vcc : std_logic;
signal XA : std_logic_vector(10 downto 0);
signal D0 : std_logic_vector(7 downto 0);
signal D1 : std_logic_vector(7 downto 0);
signal EN : std_logic;

begin

	--
	-- fixed signals
	--
	net_gnd<=(others=>'0');
	net_vcc<='1';
	--
	-- reverse address signal
	--
	XA<=A(10 downto 5)&(not A(4 downto 0));
	D<=D0 when A(11)='0' else D1;
	EN<=not CS;

	--
	-- RAM (1st half)
	--
   RAMB16_S9_inst0 : RAMB16_S9
	generic map (
		INIT => X"000", --  Value of output RAM registers at startup
		SRVAL => X"000", --  Ouput value upon SSR assertion
		WRITE_MODE => "NO_CHANGE",
		INIT_00 => X"C34A00C3E607C30E09C31809C32009C32409C33509C39308C3A108C3BD08C332",
		INIT_01 => X"0AC33604C37504C3D804C3F804C38805C3C701C308030000C33810C35803C377",
		INIT_02 => X"05C3E502C3AB02C3BE0231F010ED56CD3E07CD320A3019FE202015D3E111F0FF",
		INIT_03 => X"216B00010500EDB0C3F0FFD3E0C3000006FF21F110CDD80F3E16CD12003E7121",
		INIT_04 => X"00D8CDD509218D033EC33238102239103E04329E11CDBE02CD090011E706DFCD",
		INIT_05 => X"77053E01329D112100E8771855CD09003E2ACD120011A311CD03001A13FE0D28",
		INIT_06 => X"ECFE4A282EFE4C2848FE462832FE422826FE232886FE50287CFE4DCAA807FE53",
		INIT_07 => X"CA5E0FFE56CACB0FFE44CA290D0000000018C8CD3D01E93A9D111F3F1718A521",
		INIT_08 => X"00F07EB720A7E9FE0228A2114701DF189CCDD80438F1CD090011A009DF11F110",
		INIT_09 => X"DFCDF80438E12A06117CFE1238E1E9E3C111A311CD03001AFE1B28D3E9FDE3F1",
		INIT_0A => X"CD100438CAFDE9434845434B2053554D2045522E0D1AFE262016131AFE4C2816",
		INIT_0B => X"FE532817FE432823FE472818FE542810CDA501C3AD0011700418F511D50318F0",
		INIT_0C => X"3E0418023E02CD8F0118CF3E1D18F70E0047CDB60178D3FF3E80D3FE0E01CDB6",
		INIT_0D => X"01AFD3FEC9D5C5F51ACD8F011A13FE0D20F6F1C1D1C9DBFEE60DB9C8CD1E0020",
		INIT_0E => X"F531F010C3AD00C5D5E53E0232A01106011AFE0D283BFEC82837FECF2827FE2D",
		INIT_0F => X"2823FE2B2827FED72823FE23216C02200421840213CD1C0238D7CDC8023815CD",
		INIT_10 => X"AB024118CC3E0332A0111318C43E0118F6CDC802F5CDBE02F1C39B06C506081A",
		INIT_11 => X"BE280923232310F83713C1C923D55E2356EB7CB728093AA0113D28032918FA22",
		INIT_12 => X"A11121A01136022BD1131A47E6F0FE3028037E18051378E60F77219C02856F4E",
		INIT_13 => X"3A9E1147AF8110FDC14FAFC9434608445F0745910646330647860541EC044264",
		INIT_14 => X"0452000043CF0744F50645330646DA0547370541A50442230452000001020304",
		INIT_15 => X"06080C10182013131313C92AA1117CB7280CD5EB2104E073723E01D118063E36",
		INIT_16 => X"3207E0AF3208E0C92100E036F8237EE681200237C93A08E00F38FA3A08E00F30",
		INIT_17 => X"FA10F2AFC9F5C5E60F473E0890329E11C1F1C92173113A7211856F7E23CB16B6",
		INIT_18 => X"CB1E0FEB2A7111C9F3C5D5E5329B113EF0329C1121C0A8AFED52E500EB2107E0",
		INIT_19 => X"367436B02B73722B360A3600232336802B4E7EBA20FB79BB20F72B00000036FB",
		INIT_1A => X"363C23D14E7EBA20FB79BB20F7E1D1C1FBC9D741300D0000E52107E036802BF3",
		INIT_1B => X"5E56FB7BB2280EAF21C0A8ED523810EB3A9B11E1C911C0A83A9B11EE01E1C9F3",
		INIT_1C => X"2106E07E2F5F7E2F57FB1318EBF5C5D5E5219B117EEE01772107E036802BE55E",
		INIT_1D => X"5621C0A8192B2BEBE17372E1D1C1F1FBC9CD20097ECDC3037EC97CCDC3037D18",
		INIT_1E => X"020000F50F0F0F0FCDDA03CD1200F1CDDA03C31200010909090DE60FFE0A3802",
		INIT_1F => X"C607C630C9D630D8FE0A3FD0D607FE103FD8FE0AC90000000018EA7F20504C41",
		INIT_20 => X"590D7F205245434F52442E0D00000000D5CD1F04380767CD1F0438016FD1C9C5",
		INIT_21 => X"1A13CDF903380D0F0F0F0F4F1A13CDF9033801B1C1C9F3D5C5E516D71ECC21F0",
		INIT_22 => X"10018000CD1A07CD9F0638187BFECC200DCD0900D5116704DF11F110DFD1CD7A",
		INIT_23 => X"07CD8A04C3540557524954494E47200D0109090B0DF3D5C5E516D71E53ED4B02",
		INIT_24 => X"112A041178B1284A18BAD5C5E516023EF83200E07ECD67073A01E0E681C2A504",
		INIT_25 => X"3E0237182D230B78B1C294042A97117CCD67077DCD6707CD1A0A15C2C204B7C3",
		INIT_26 => X"D2040600CD010A05C2C404E1C1C5E5C39404E1C1D1C92F4EF3D5C5E516D21ECC",
		INIT_27 => X"01800021F010CD9F06DA7205CD5B06DA7205CD0E05C35405F3D5C5E516D21E53",
		INIT_28 => X"ED4B02112A041178B1CA540518D8D5C5E526020101E01102E0CD01063854CD4A",
		INIT_29 => X"0A1AE620CA190554210000229711E1C1C5E5CD2406383B77230B78B120F42A97",
		INIT_2A => X"11CD2406382C5FCD24063826BD20167BBC2012AFE1C1D1CD0007F53A9C11FEF0",
		INIT_2B => X"2001FBF1C915280662CDE20F18A53E0118023E023718DDD5115203F7D1C9CDFF",
		INIT_2C => X"09CDCA08FEF0C900F3D5C5E5ED4B02112A041116D21E5378B128B9CD1A07CD9F",
		INIT_2D => X"0638CFCD5B0638CACDAD0518A7D5C5E526020101E01102E0CD0106DA7205CD4A",
		INIT_2E => X"0A1AE620CAB80554E1C1C5E5CD240638A1BE209A230B78B120F22A9911CD2406",
		INIT_2F => X"BC208BCD2406BD208515CA53056218C2F53A8E11CDB10F77F1C9CD0900CDBA03",
		INIT_30 => X"C93EF83200E0000AE681200237C91AE62020F40AE681200237C91AE62028F4C9",
		INIT_31 => X"00000000C5D5E52100080101E01102E0CD0106DA5406CD4A0A1AE620CA4906E5",
		INIT_32 => X"2A971123229711E1377D176F25C23006CD01067DE1D1C1C9000000CDE20FC5D5",
		INIT_33 => X"E52128287BFECC28032114142295110101E01102E02A9511CD0106381ECD4A0A",
		INIT_34 => X"1AE62028F02520F0CD0106380ECD4A0A1AE62020E02D20F0CD0106E1D1C1C9C5",
		INIT_35 => X"D5E5060A3A02E0E610280E06FFCD9609180218EB10F7AF18E23E062103E0773C",
		INIT_36 => X"7710E1CD09007AFED7280511FB031807110204DF11FD03DF3A02E0E61020CCCD",
		INIT_37 => X"320A20F43718D02A2A20204D4F4E49544F5220315A2D3031334120202A2A0D00",
		INIT_38 => X"F5C5D5060A3A02E0E610280B3E063203E03C3203E010EEC3E60EC5D5E5110000",
		INIT_39 => X"78B1200BEB229711229911E1D1C1C97EC506080730011310FAC1230B18E22103",
		INIT_3A => X"E0368A36073605C900000000000000000000000000000000003E153DC25B07C9",
		INIT_3B => X"3E133DC26207C9C50608CD1A0A07DC1A0AD4010A05C26D07C1C9C5D57B01F055",
		INIT_3C => X"112828FECCCA8E0701F82A111414CD010A0B78B120F8CD1A0A1520FACD010A1D",
		INIT_3D => X"20FACD1A0AD1C1C9CD3D01CDFA05CDB103CD2009CD2F01CD1004381BCDA60213",
		INIT_3E => X"CD1F0438E6BE20E3131AFE0D2806CD1F0438D8772318D4606918D028484C29F1",
		INIT_3F => X"9E5355422028F5C5E5D5CDB309F5473A9D110FD4770578217011E6F0FEC0D178",

		INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")

	port map (
		DO => D0,				-- 8-bit Data Output
		DOP => open,			-- 1-bit parity Output
		ADDR => XA,	-- 11-bit Address Input
		CLK => CLK,			-- Clock
		DI => net_gnd(7 downto 0),		-- 8-bit Data Input
		DIP => net_gnd(0 downto 0),		-- 1-bit parity Input
		EN => EN,		-- RAM Enable Input
		SSR => net_gnd(0),		-- Synchronous Set/Reset Input
		WE => net_gnd(0)		-- Write Enable Input
	);

	--
	-- RAM (2nd half)
	--
   RAMB16_S9_inst1 : RAMB16_S9
	generic map (
		INIT => X"000", --  Value of output RAM registers at startup
		SRVAL => X"000", --  Ouput value upon SSR assertion
		WRITE_MODE => "NO_CHANGE",
		INIT_00 => X"2016FECD2855FECBCA2208FECF2809FEC7300ACB1B783005CDB50D18CDCDDC0D",
		INIT_01 => X"18C8E1E5361B23360D18530F30371833CD9609CD500AC9000000000000000000",
		INIT_02 => X"000000000000000000000000000000000000000000000000000000CDF3020628",
		INIT_03 => X"30C92506502E00CDB40FD1D57ECDCE0B12231310F7EB360D2B7EFE2028F8CD0E",
		INIT_04 => X"09D1E1C1F1C900000000000000000000000000F5C5D51AFE0D280CCD35091318",
		INIT_05 => X"F5F5C5D51AFE0DCAE60ECDB90BCD6C091318F1112A0C18423ECBB71819CDCA08",
		INIT_06 => X"D6F0C8C6F0C3CE0B0000C5D5E5CD3008780738063EF0E1D1C1C911EA0B78FE88",
		INIT_07 => X"28D6260069CB6F200E3A70110FDAFE0878171738BE180311AA0C197E18D8CB70",
		INIT_08 => X"280711E90C193718F2116A0C18ECAF3294113ECD184300003A9411B7C818EF00",
		INIT_09 => X"3E201811CD0C003A9411B7C8D60A38F420FA000000FE0D28D5C54F47CD460978",
		INIT_0A => X"C1C94F4B210D79CDB90B4FFEF0C8E6F0FEC0792017FEC73013CDDC0DFEC3280F",
		INIT_0B => X"FEC52803FEC6C0AF329411C9CDB50D3A94113CFE5038F1D65018ED3A8E11186F",
		INIT_0C => X"CB6F2802B7C93E20B737C946494C454E414D453F200DC50615CD4A0A10FBC1C9",
		INIT_0D => X"4C4F4144494E47200D3E593DC2AB09C9000000E5CD920BCD7E0520FBCD7E0528",
		INIT_0E => X"FB67CD9609CDCA08F5BCE120EFE5F1CDF005E1C9AF010008D55772230B78B120",
		INIT_0F => X"F9D1C9F5E53A02E00707388F3A9211CDB10F77E1F1C900000000000000000018",
		INIT_10 => X"E2F53E033203E0CD5907CD59073E023203E0CD5907CD5907F1C9F53E033203E0",
		INIT_11 => X"CDA9093E023203E0CDA909F1C900000000003EF83200E0003A01E0B71FDA8009",
		INIT_12 => X"171730043E4037C9AFC93E3FC3620700D5E5AF06F857CD320A20041688181430",
		INIT_13 => X"05571802CBFA05783200E0FEEF2008FEF828F342E1D1C93A01E02FB728E85F26",
		INIT_14 => X"0878E60F0707074F7B250F30FC7C814F18D2F0F0F0F3F0F5F0F0F0F0F0F0F0F0",
		INIT_15 => X"F0F0F0C1C2C3C4C5C6F0F0F0F0F0F0F0F0F0006162636465666768696B6A2F2A",
		INIT_16 => X"2E2D202122232425262728294F2C512B5749550102030405060708090A0B0C0D",
		INIT_17 => X"0E0F101112131415161718191A5259545045C7C8C9CACBCCCDCECFDFE7E8E5E9",
		INIT_18 => X"ECEDD0D1D2D3D4D5D6D7D8D9DADBDCDDDEC080BD9DB1B5B9B49EB2B6BABE9FB3",
		INIT_19 => X"B7BBBFA385A4A5A69487889C82988492908391819A97939589A1AF8B8696A2AB",
		INIT_1A => X"AA8A8EB0AD8DA7A8A98F8CAEAC9BA099BCB8403B3A703C715A3D43563F1E4A1C",
		INIT_1B => X"5D3E5C1F5F5E377B7F367A7E334B4C1D6C5B7841353474303875394D6F6E3277",
		INIT_1C => X"767273477C53314E6D48467D441B5879426021921136EF3A70110F38030F3002",
		INIT_1D => X"36FF7EF5CDB10F7E328E11F177AF2100E0772F77C9364318E9C5E521920A4F06",
		INIT_1E => X"00097E181B56312E30410D000000C5E5D521920A545D010001EDB128063EF0D1",
		INIT_1F => X"E1C1C9B72BED527D18F5BFCA58C9F02C4FCD191A555254F0F0F0111213141516",
		INIT_20 => X"1718090A0B0C0D0E0F100102030405060708212223242526272859502A002029",
		INIT_21 => X"2F2EC8C7C2C1C3C4492DBFCA1BC9F06A6BCD999AA4BC40F0F0F0919293949596",
		INIT_22 => X"9798898A8B8C8D8E8F908182838485868788616263646566676880A52B006069",
		INIT_23 => X"5157C6C5C2C1C3C45A45BFF0E5C9F042B6CD7576B2D84EF0F0F03C30447179DA",
		INIT_24 => X"386D7D5C5BB41C32B0D6536FDE47344A4B72373E7F7B3A5E1FBDD49ED2009CA1",
		INIT_25 => X"CAB8C8C7C2C1C3C4BADBF0F0F0F0F0F0F0F0F05AF0F0F0F0F0F0C1C2C3C4C5C6",
		INIT_26 => X"F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0",
		INIT_27 => X"F0F0F0F0F0F0F0F0F0BFF0CFC9F0B54DCD3577D7B3B7F0F0F07C70413139A678",
		INIT_28 => X"DD3D5D6C561D33D5B1466ED94874434C733F367E3B7A1E5FA2D39FD1009DA3D0",
		INIT_29 => X"B9C6C5C2C1C3C4BBBECD3D01CDA602E5CD1004D13852EB06080E17CDFA05CDB1",
		INIT_2A => X"0323F53A711181327111F1FE2030023E2ECDB90BCD6C093A71110C913271110D",
		INIT_2B => X"0D0DE5ED52E1281D3EF83200E0003A01E0FEFE2003CDA60D10C4CDCA08B728FA",
		INIT_2C => X"CD320A20B2C3AD0021A0001918A8000000000000000000000000000000000000",
		INIT_2D => X"000000000000F53A02E00730FA3A02E00738FAF1C9F5C5D5E5CDB10F772A7111",
		INIT_2E => X"7DFE27200BCDF3023806EB36012336003EC3180C3A7011FE013ECAC9F5C5D5E5",
		INIT_2F => X"47E6F0FEC0201BA8074F060021AA0E095E23562A7111EBE9EB7CFE1828252422",
		INIT_30 => X"7111C3E50EEB7CB728F82518F2EB7DFE2730032C18E92E00247CFE1938E12618",
		INIT_31 => X"2271111848EB7DB728032D18D22E2725F20B0E260022711118C8217311061BCD",
		INIT_32 => X"D80F2100D0CDD4093E71CDD50921000018AD0000000000000000CDF3020F30B6",
		INIT_33 => X"2E0024FE18280324189522711101C0031100D02128D0C5EDB0C1D51100D82128",
		INIT_34 => X"D8EDB00628EB3E71CDDD0FE10628CDD80F011A00117311217411EDB036003A73",
		INIT_35 => X"11B728412172113518C36D0EF80D050E0D0E250E4D0E3A0EF80E380FE10EEE0E",
		INIT_36 => X"E50EE50E5A0EE50EE50ECBDC7E23772BCB9CEDA879B020F2EB3600CBDC367118",
		INIT_37 => X"04AF327011E1D1C1F1C900000000CDD40DCAB90D3E0118EAEB7CB528E87DB720",
		INIT_38 => X"0DCDF3023808CDB10F2B36001825CDF3020F3E283001079547CDB10F7E2B7723",
		INIT_39 => X"CBDC7E2B77CB9C232310F12B3600CBDC2171003EC4C3E00DCDF3020F2E277D30",
		INIT_3A => X"0124CDB40FE52A711130023E4F9506004FD128911AB7208D626B2BC3CA0ECD3D",
		INIT_3B => X"01220411444DCDA602CD3D01ED4223220211CDA602CD3D01220611CD0900118B",
		INIT_3C => X"09DFCD2F01CDA602CDA60221F110131A7723FE0D20F83E0132F010CD3604DA07",
		INIT_3D => X"01CD7504DA0701CD0900114209DFC3AD002A7111F5C5D5E5C111280021D8CF19",
		INIT_3E => X"05F2BF0F060009D1C1F1C9CD8805DA0701114209DFC3AD00AF18023EFF772310",
		INIT_3F => X"FCC9C5D5E50101E01102E02664CD0106380BCD4A0A1AE62020F12520F0C39B06",

		INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")

	port map (
		DO => D1,				-- 8-bit Data Output
		DOP => open,			-- 1-bit parity Output
		ADDR => XA,	-- 11-bit Address Input
		CLK => CLK,			-- Clock
		DI => net_gnd(7 downto 0),		-- 8-bit Data Input
		DIP => net_gnd(0 downto 0),		-- 1-bit parity Input
		EN => EN,		-- RAM Enable Input
		SSR => net_gnd(0),		-- Synchronous Set/Reset Input
		WE => net_gnd(0)		-- Write Enable Input
	);

end Behavioral;

