--
-- mom.vhd
--
-- MONITOR 1Z-009A/MZ NEW-MONITOR module
-- for MZ-700 on FPGA
--
-- Nibbles Lab. 2005
--

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

--  Uncomment the following lines to use the declarations that are
--  provided for instantiating Xilinx primitive components.
library UNISIM;
use UNISIM.VComponents.all;

entity mrom is
    Port ( A : in std_logic_vector(11 downto 0);
           CS : in std_logic;
           D : out std_logic_vector(7 downto 0);
		 CLK : in std_logic);
end mrom;

architecture Behavioral of mrom is

--
-- signals
--
signal net_gnd : std_logic_vector(7 downto 0);
signal net_vcc : std_logic;
signal XA : std_logic_vector(10 downto 0);
signal D0 : std_logic_vector(7 downto 0);
signal D1 : std_logic_vector(7 downto 0);
signal EN : std_logic;

begin

	--
	-- fixed signals
	--
	net_gnd<=(others=>'0');
	net_vcc<='1';
	--
	-- reverse address signal
	--
	XA<=A(10 downto 5)&(not A(4 downto 0));
	D<=D0 when A(11)='0' else D1;
	EN<=not CS;

	--
	-- RAM (1st half)
	--
   RAMB16_S9_inst0 : RAMB16_S9
	generic map (
		INIT => X"000", --  Value of output RAM registers at startup
		SRVAL => X"000", --  Ouput value upon SSR assertion
		WRITE_MODE => "NO_CHANGE",
		INIT_00 => X"C300E8C3E607C30E09C31809C32009C37F00C33509C38109C39909C3BD08C332",
--		INIT_00 => X"C34A00C3E607C30E09C31809C32009C37F00C33509C38109C39909C3BD08C332",
		INIT_01 => X"0AC33604C37504C3D804C3F804C38805C3C701C308030000C33810C35803C3E5",
		INIT_02 => X"02C3FA02C3AB02C3BE0231F010ED56CDC90F3E16D7063C217011CDD80F219203",
		INIT_03 => X"3EC3323810223910210405229E11CDBE02114101DFCDC00A180811F1101896C3",
		INIT_04 => X"260931F010118200D5CD09003E2AD711A311CD03001AFE2AC2540C131AFE47CA",
		INIT_05 => X"5901FE23CA1202FE4DCA0F0CFE53CA820CFE26CA0E0EFE4C281F00000000FE52",
		INIT_06 => X"CAAA01FE50CA1202C39B0ACDE800CD2D00380A11C401CFDFC9CDE800EFDA6701",
		INIT_07 => X"2A06117CFE12D8E9CD27003895CF113801DF18861100D00E1906281ACDCE0BCD",
		INIT_08 => X"0F011310F63E0DCD0F010D20ECC9D5F5DBFEE60DB72807CD1E00287718F2F1D3",
		INIT_09 => X"FF3E80D3FEDBFEE60DFE0120F8AFD3FEC9464F554E44200D4C4F2E200DC34901",
		INIT_0A => X"00204D5A903730300DD3E111F0FFD5212E07010500EDB0C900131AFE4F200413",
		INIT_0B => X"131313CDC00CE9FE02C8CF11B501DFC93EFF329D11C9AF18F92100F07EB7C0E9",
		INIT_0C => X"C5D5E51ABE200B052808FE0D2804132318F1E1D1C1C9F5C3AD0D3EFFD3E0C911",
		INIT_0D => X"3101DF11F110DFC3E30FCDE800CDE30FEFC3D1000043450D36FF3A7011B72002",
		INIT_0E => X"36EFAFC94F4B0DC5D5E53E0232A01106011AFE0D2802FEC8282EFECF281EFED7",
		INIT_0F => X"2822FE2321710220032E8913CD1C0238E0CDC8023815CDAB024118D53E0332A0",
		INIT_10 => X"111318CD3E0118F6CDC802F5CDBE02F1188013CD1F04D8CD0F0118F6C506081A",
		INIT_11 => X"BE280923232310F83713C1C923D55E2356EB7CB728093AA0113D28032918FA22",
		INIT_12 => X"A1113E0232A011D1131A47E6F0FE3028053A9F1118071378E60F329F114F0600",
		INIT_13 => X"21A102094E3A9E1147AF8110FDC14FAFC943770744A70645ED0546980547FC04",
		INIT_14 => X"41710442F503520000430C0744470645980546480547B40441310442BB035200",
		INIT_15 => X"000102030406080C1018202AA1117CB7280CD5EB2104E073723E01D118063E36",
		INIT_16 => X"3207E0AF3208E0C92100E036F8237EE680200237C93A08E00F38FA3A08E00F30",
		INIT_17 => X"FA10F2AFC9C5E5217104CDAE020632AFCD5B0710FAE1C1C3BE02F5C5E60F473E",
		INIT_18 => X"0890329E11C1F1C9F3C5D5E5329B113EF0329C1121C0A8AFED52E523EB3E7432",
		INIT_19 => X"07E03EB03207E02106E073722B360A36003E803207E0234E7EBA20FB79BB20F7",
		INIT_1A => X"2B0000003612367A23D14E7EBA20FB79BB20F7E1D1C1FBC9E53E803207E02106",
		INIT_1B => X"E0F35E56FB7BB2CA7903AF21C0A8ED52DA8303EB3A9B11E1C911C0A83A9B11EE",
		INIT_1C => X"01E1C9F32106E07E2F5F7E2F57FB13C37C03F5C5D5E53A9B11EE01329B113E80",
		INIT_1D => X"3207E02106E05E5621C0A8192B2BEB2106E07372E1D1C1F1FBC97CCDC3037DCD",
		INIT_1E => X"C303C9F5E6F00F0F0F0FCDDA03CD1200F1E60FCDDA03D73E20C9D5E521E903E6",
		INIT_1F => X"0F5F1600197EE1D1C930313233343536373839414243444546C5E501001021E9",
		INIT_20 => X"03BE2003791806230C0520F537E1C1C9D5CD1F04380767CD1F0438016FD1C9C5",
		INIT_21 => X"1A13C3F106380D070707074F1A13CDF9033801B1C1C9F3D5C5E516D71ECC21F0",
		INIT_22 => X"10018000CD3307CDB206DA63057BFECC2011CD0900D5116C04CD150011F110CD",
		INIT_23 => X"1500D1CDB807CD8D04C3630557524954494E47200DF3D5C5E516D71E532A0211",
		INIT_24 => X"E5C12A041178B1CAD404C34404D5C5E53A3710573EF83200E07ECDA5073A01E0",
		INIT_25 => X"E608200337182D230B78B1C299042A97117CCDA5077DCDA507CD800715C2C404",
		INIT_26 => X"B7C3D4040600CD670705C2C604E1C1C5E5C39904E1C1D1C9F3D5C5E516D21ECC",
		INIT_27 => X"01800021F010CDB206DA8205CD5E06DA8205CD1005C36305F3D5C5E516D21E53",
		INIT_28 => X"2A0211E5C12A041178B1CA6305C3E604D5C5E52A36100101E01102E0CD010638",
		INIT_29 => X"61CD55061AE62028F354210000229711E1C1C5E5CD2406384977230B78B120F4",
		INIT_2A => X"2A9711CD2406383A5FCD24063834BD20237BBC201F180B3E01323710C93E0218",
		INIT_2B => X"F800AFE1C1D1CD0007F53A9C11FEF02001FBF1C915CA7C0562C316053E0137C3",
		INIT_2C => X"63053E0237C36305F3D5C5E52A0211E5C12A041116D21E5378B1CA6305CD3307",
		INIT_2D => X"CDB206DA8205CD5E06DA8205CDB205C36305D5C5E52A36100101E01102E0CD01",
		INIT_2E => X"0638BFCD55061AE62028F354E1C1C5E5CD240638ADBE20A4230B78B120F22A99",
		INIT_2F => X"11CD2406BC2095CD2406BD208F15CA620562C3B8057806C0803002D64047C33A",
		INIT_30 => X"083EF93200E0000AE604C20F0637C91AE620C207060AE608C21D0637C91AE620",
		INIT_31 => X"CA1506C9C5D5E52100080101E01102E0CD0106381CCD55061AE620280AE52A97",
		INIT_32 => X"1123229711E1377D176F2520E3CD01067DE1D1C1C93A35103D20FD2000C9C5D5",
		INIT_33 => X"E52128287BFECC28032114142295110101E01102E02A9511CD0106381ECD5506",
		INIT_34 => X"1AE62028F02520F0CD0106380ECD55061AE62020E02D20F0CD0106E1D1C1C9C2",
		INIT_35 => X"F5053E282A71119547CDB10FCDD80FC3EE07C5D5E50E0A3A02E0E6102805AFE1",
		INIT_36 => X"D1C1C93E062103E0773C770D20E9CF7AFED72806112207DF1808112907DF1124",
		INIT_37 => X"07DF3A02E0E61020D5CD440A20F43718CEFE2F2806CDF903C325041A13C33404",
		INIT_38 => X"F5C5D5060A3A02E0E6102004D1C1F1C93E063203E03E073203E005C20507D1C1",
		INIT_39 => X"F1C97F20504C41590D7F5245430DD3E0C30000C5D5E511000078B1200BEB2297",
		INIT_3A => X"11229911E1D1C1C97EE52608073001132520F9E1230B18E13A36103D20FDC93A",
		INIT_3B => X"370018F4000000F53E033203E0CD5F073E023203E0CD5F07F1C908C3E4090000",
		INIT_3C => X"F53E033203E0CD5F07CD5F073E023203E0CD5F07CD6207F1C93E003234102144",
		INIT_3D => X"2E223510C9C50608CD800707DC8007D4670705C2AB07C1C9C5D57B01F82A1128",
		INIT_3E => X"28FECCCACC0701BE0A111414CD67070B78B120F8CD80071520FACD67071D20FA",
		INIT_3F => X"CD8007D1C1C9F5C5E5D5AF329311CDB309473A9D11B7CC6D0C78E6F0FEC02037",
		INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
	port map (
		DO => D0,				-- 8-bit Data Output
		DOP => open,			-- 1-bit parity Output
		ADDR => XA,	-- 11-bit Address Input
		CLK => CLK,			-- Clock
		DI => net_gnd(7 downto 0),		-- 8-bit Data Input
		DIP => net_gnd(0 downto 0),		-- 1-bit parity Input
		EN => EN,		-- RAM Enable Input
		SSR => net_gnd(0),		-- Synchronous Set/Reset Input
		WE => net_gnd(0)		-- Write Enable Input
	);

	--
	-- RAM (2nd half)
	--
   RAMB16_S9_inst1 : RAMB16_S9
	generic map (
		INIT => X"000", --  Value of output RAM registers at startup
		SRVAL => X"000", --  Ouput value upon SSR assertion
		WRITE_MODE => "NO_CHANGE",
		INIT_00 => X"78FECD2856FEC9281DFECA2814FECBCAB308FEC8280BFEC728073A9311B7201C",
		INIT_01 => X"78CDDC0D18C8217011AFBE20013C77D6062F3203E018B7CD440A286A78CDA60D",
		INIT_02 => X"CDB50DFE6220A72193117E2F77189FFE10CA420FFED5FE05C39F062A71115C16",
		INIT_03 => X"0021731119EB1AB70128002A7111C27A08131AB7CA7D08C37B08250E502E00CD",
		INIT_04 => X"B40FD1D5C5CDA60DEDB0C1E1E5417ECDCE0B772310F8360D2B7EFE2028F8CD06",
		INIT_05 => X"00D1E1C1F1C978FE12CAF60DFE49CA290E189CE1E5361B23360D18E200CDCA08",
		INIT_06 => X"FEF02002AFC9CDCE0BC9C5D5E5CD500A780738063EF0E1D1C1C907D2EC080600",
		INIT_07 => X"2108000911C90A197EC3D6083A7011B7C2FD08060021C90A097EC3D60879E6F0",
		INIT_08 => X"0F4779E60F80C6A06F2600C3E408AF3294113ECDCDDC0DC93A9411B7C8C30600",
		INIT_09 => X"3E20CD3509C9CD0C003A9411B7C8D60A38F420FAC9FE0DCA0E09C54F47CD9601",
		INIT_0A => X"CD460979C1C979CDB90B4FE6F0FEF0C8FEC079C27009FEC7D27009CDDC0DFEC3",
		INIT_0B => X"CA7309FEC5CA6B09FEC6C0AF329411C9CDB50D3A94113CFE503802D650329411",
		INIT_0C => X"C9F5C5D50605CD96011AFE0DCADF0F4FCD46091310F3C38409F5C5D50605CD96",
		INIT_0D => X"011AFE0DCADF0FCDB90BCD70091310F1C39C09C5D5E5CDB10FCDA60D7E328E11",
		INIT_0E => X"228F11219211CDB8013200E03291112F3200E01614CDFF09CD500A7807DAE60B",
		INIT_0F => X"15C2D509CDFF09CDCA08FEF0CA7A07F5CDA60D3A8E112A8F1177F1E1D1C1C9F5",
		INIT_10 => X"E53A02E00707DA250A3A91110FDA220A3A92112A8F11CDA60D773A9111EE0132",
		INIT_11 => X"9111E1F1C93A91110FD2220A3A8E11C3130A3EF83200E0003A01E02FE621C244",
		INIT_12 => X"0AC601C93EF83200E0003A01E0E680C9D5E506FA160005783200E0FEEF200442",
		INIT_13 => X"E1D1C9FEF8281F3A01E02FB728E85FCBFA78E60F070707074F3E083D2804CB03",
		INIT_14 => X"30F9814F18D03A01E02F5FE6212802CBF27BE6DE28C018D6CD3E00FE56CACB00",
		INIT_15 => X"FE43C0131AFE41CA9E07FE31CA5705FE32CA5D05FE42C2B80C212215223510C9",
		INIT_16 => X"CD9907CD5D05C37601CD4F2CF0C92BF0CACD1B39F0C93EF0CAF0F0F06968551A",
		INIT_17 => X"19F0F0F04A366D5A3D181716151413121153734670715D3372100F0E0D0C0B0A",
		INIT_18 => X"0976774356785E1E3C08070605040302015F1F1D321C44415C28272625242322",
		INIT_19 => X"2152676665646362612E2F2920002A6A6B5751546000DDDE592D49C4C3C1C2C7",
		INIT_1A => X"C84540C4C3C1C2C5C6F0C7F0C3CDF0F0F0F0C8F0C4CDF0F0CBC500C1CBF03C3E",
		INIT_1B => X"DCC600C2F0F07C7ED8CDBC8DF0C999F0CAF0F0F0B8B4A091868187979682849C",
		INIT_1C => X"94AAAB8F8CADB08EA28A839088929A9398A18995A6A5A485A3ACAEAF8B00A7A8",
		INIT_1D => X"A99BBFC4C3C1C2C7C8F0C7F0C3CDF0BDBFC500C1F0F0BCBEDBC5E5FE17381C21",
		INIT_1E => X"C60C01E000EDB1201A3EDF91180AC5E521C60C4F0600097EE1C1C9FE113804C6",
		INIT_1F => X"B018F5AF18F23A3410B7C2D3097908B9CAE0090604CDCA08E63F57CDFF09CDCA",
		INIT_20 => X"08E63FBAC2E7090B78B1CAE40918EC13CD10040610CD300CCDCA08B72805FECB",
		INIT_21 => X"C810F2CDB309FECD28E9B7C0060118E5C5CDBA030608C5E5AFD77ECDC30323AF",
		INIT_22 => X"D710F7D7E1C17ECDB90BCDB50D2310F6C1C30600CDC00C1EA8CD1F0438057713",
		INIT_23 => X"2318F63EA9BBD0CDBA03C38E00C5E52A36107DFE1038032E5024CDAE020607C3",
		INIT_24 => X"EF02131AFE53CA7001FE47CA7601CDC00C220411E51EAACD1004D1ED52232202",
		INIT_25 => X"1111AF11CDC00C22061111F11021B411011000EDB03E0D12CD9F01E7D22400C9",
		INIT_26 => X"CD1004D0D1C9204142434445464748494A4B4C4D4E4F50515253545556575859",
		INIT_27 => X"5AFBCDDDCBD1303132333435363738392D3D3B2F2E2CE5F4ECDAE3E2D7D4E6E8",
		INIT_28 => X"C2C1C4C7CFCA20E1FEC8FA5FF8F1F73FCCDBDCE9F53A5E3C5BF35D40C93EFC5C",
		INIT_29 => X"C6DFD0CED3D2FF2122232425262728292B2ADEF6EBEAC3C5EFF0E4E7EEEDE0FD",
		INIT_2A => X"D8D5F2F9D9D620A19A9F9C92AA9798A6AFA9B8B3B0B79EA09DA496A5ABA39BBD",
		INIT_2B => X"A2BB9982878CBCA7AC91939495B4B5B6AEADBAB2B9A8B183888D8684898EBF85",
		INIT_2C => X"8A8FBE818B907F11121314151660616263646566676870711173747576777879",
		INIT_2D => X"7A7B7C7D7E69F53A02E00730FA3A02E00738FAF1C9F5C5D5E547CDB10F702A71",
		INIT_2E => X"117DFE27C2900E5C1600217311197EB7C2900E233601233600C3900EF5C5D5E5",
		INIT_2F => X"47E6F0FEC0207FA8FE0DCA8B0FFE0B3075260E6F6EE92134107E2F77C3EE0700",
		INIT_30 => X"32748490AEBFC5F80BE1F2C3490F11A311D5211B0E010C00EDB0C92102E0CB9E",
		INIT_31 => X"CBC6CB86C38009DF00219D1118CB00C37D08CD9601AF3203E001C0031100D021",
		INIT_32 => X"28D0EDB0EB0628CDD80F011A00117311217411EDB036003A7311B7C26A0ECD96",
		INIT_33 => X"013E013203E0C3DE0F002A711125227111C3390E2A71117CFE18CA320E242271",
		INIT_34 => X"11C3DE0F2A71117CB7CADE0F25C37E0E2A71117DFE27D29D0E2CC37E0E2E0024",
		INIT_35 => X"7CFE19DA7E0E2618227111C3320E2A71117DB728042DC37E0E2E2725F27E0E21",
		INIT_36 => X"0000C37E0ECDA60D0E192100D00628CDD80F0DC2CD0E217311061BCDD80FC3BF",
		INIT_37 => X"0E217011AFBE18013C77D6062F3203E0188F217011AF18F02A71117CB5CADE0F",
		INIT_38 => X"7DB720165C1600217311197EB7200BCDB10FCDA60D2B360018942A71115C1C16",
		INIT_39 => X"00217311197E47B73E2828023E502A7111954F0600CDB10FE5D11BCDA60DEDB0",
		INIT_3A => X"18D3CDF400C3EE07002A71115C1C1600217311197EB70E002A71112E27280224",
		INIT_3B => X"0CCDB40F7EB7C2DE0FE52A71113E27954779B728043E288047D1D5E12BCDA60D",
		INIT_3C => X"7E1236002B1B10F8C3DE0F2A71115C1C1600217311197EB72A7111CA9D0E2E00",
		INIT_3D => X"7CFE1728052424C37E0E24227111C3320E2A7111C5D5E5C111280021D8CF1905",
		INIT_3E => X"F2BE0F060009D1C1C92103E0368A360736053E013203E0C9AF772310FCC9E1D1",
		INIT_3F => X"C1F1C93E3AD72A0411CDBA03EB2A0211192BCDF80F2A06113E2DD7CDBA03AFC9",
		INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
	port map (
		DO => D1,				-- 8-bit Data Output
		DOP => open,			-- 1-bit parity Output
		ADDR => XA,	-- 11-bit Address Input
		CLK => CLK,			-- Clock
		DI => net_gnd(7 downto 0),		-- 8-bit Data Input
		DIP => net_gnd(0 downto 0),		-- 1-bit parity Input
		EN => EN,		-- RAM Enable Input
		SSR => net_gnd(0),		-- Synchronous Set/Reset Input
		WE => net_gnd(0)		-- Write Enable Input
	);

end Behavioral;
