--
-- cgrom.vhd
--
-- MZ-700 CG-ROM pattern module
-- for MZ-700 on FPGA
--
-- Nibbles Lab. 2005
--

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

--  Uncomment the following lines to use the declarations that are
--  provided for instantiating Xilinx primitive components.
library UNISIM;
use UNISIM.VComponents.all;

entity cgrom is
    Port ( ROMA : in std_logic_vector(10 downto 0);
           CSEL : in std_logic;
           ROMD : out std_logic_vector(7 downto 0);
		 PCGSW : in std_logic;
		 CSPCG : in std_logic;
		 WR : in std_logic;
           RAMA : in std_logic_vector(1 downto 0);
           RAMD : in std_logic_vector(7 downto 0);
		 MCLK : in std_logic;
		 DCLK : in std_logic);
end cgrom;

architecture Behavioral of cgrom is

--
-- CG-ROM
--
signal net_gnd : std_logic_vector(7 downto 0);
signal net_vcc : std_logic;
signal XA : std_logic_vector(10 downto 0);
signal D0 : std_logic_vector(7 downto 0);
signal D1 : std_logic_vector(7 downto 0);
signal CPYD0 : std_logic_vector(7 downto 0);
signal CPYD1 : std_logic_vector(7 downto 0);
--
-- PCG
--
signal EXA : std_logic_vector(10 downto 0);
signal D2 : std_logic_vector(7 downto 0);
signal CPYA : std_logic_vector(10 downto 0);
signal PCGA : std_logic_vector(10 downto 0);
signal TMPA : std_logic_vector(2 downto 0);
signal BUFD : std_logic_vector(7 downto 0);
signal PCGD : std_logic_vector(7 downto 0);
signal PCGWP : std_logic;
signal PCGDSEL : std_logic;
signal TMPDSEL : std_logic;

begin

	--
	-- fixed signals
	--
	net_gnd<=(others=>'0');
	net_vcc<='1';
	--
	-- reverse address signal
	--
	XA<=ROMA(10 downto 5)&(not ROMA(4 downto 0));
	EXA<=CSEL&XA(9 downto 0);

	--
	-- Font select
	--
	process( CSEL, XA(10), PCGSW, D0, D1, D2 ) begin
		if( CSEL='0' ) then
			if( PCGSW='0' ) then
				ROMD<=D0;
			else
				if( XA(10)='0' ) then
					ROMD<=D0;
				else
					ROMD<=D2;
				end if;
			end if;
		else
			if( PCGSW='0' ) then
				ROMD<=D1;
			else
				if( XA(10)='0' ) then
					ROMD<=D1;
				else
					ROMD<=D2;
				end if;
			end if;
		end if;
	end process;

	--
	-- Access Registers
	--
	process( MCLK ) begin
		if( MCLK'event and MCLK='1' ) then
			PCGA(10 downto 8)<=TMPA;
			PCGDSEL<=TMPDSEL;
			if( CSPCG='0' and WR='0' ) then
				if( RAMA="00" ) then
					BUFD<=RAMD;
				elsif( RAMA="01" ) then
					PCGA(7 downto 0)<=RAMD(7 downto 5)&(not RAMD(4 downto 0));
				elsif( RAMA="10" ) then
					TMPA<=RAMD(2 downto 0);
					PCGWP<=not RAMD(4);
					TMPDSEL<=RAMD(5);
				end if;
			end if;
		end if;
	end process;
	CPYA<='1'&TMPA(1 downto 0)&PCGA(7 downto 0);
	PCGD<=BUFD when PCGDSEL='0' else
		 CPYD0 when PCGDSEL='1' and PCGA(10)='0' else
		 CPYD1;

	--
	-- RAM (CG data included:normal)
	--
   RAMB16_S9_S9_inst0 : RAMB16_S9_S9
	generic map (
      INIT_A => X"000", --  Value of output RAM registers on Port A at startup
      INIT_B => X"000", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"000", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"000", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "READ_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "READ_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
		INIT_00 => X"00000000000000003C42427E424242007C22223C22227C003C42404040423C00",
		INIT_01 => X"7C22222222227C007E40407840407E007E404078404040003C42404E42423C00",
		INIT_02 => X"4242427E424242001C08080808081C000E040404044438004244487048444200",
		INIT_03 => X"4040404040407E0042665A5A424242004262524A464242001824424242241800",
		INIT_04 => X"7C42427C40404000182442424A241A007C42427C484442003C42403C02423C00",
		INIT_05 => X"3E080808080808004242424242423C0042424224241818004242425A5A664200",
		INIT_06 => X"42422418244242002222221C080808007E02041820407E000C12103810103E00",
		INIT_07 => X"080808080F00000008080808F8000000080808080F08080808080808FF000000",
		INIT_08 => X"3C42465A62423C000818280808083E003C42020C30407E003C42023C02423C00",
		INIT_09 => X"404044447E0404007E407C0202423C003C40407C42423C007E42040810101000",
		INIT_0A => X"3C42423C42423C003C42423E02423C000000007E0000000000007E007E000000",
		INIT_0B => X"0000080000080810000204081020400000000000001818000000000000181830",
		INIT_0C => X"00FF000000000000404040404040404080808080808080FF01010101010101FF",
		INIT_0D => X"000000FF000000001010101010101010FFFF000000000000C0C0C0C0C0C0C0C0",
		INIT_0E => X"0000000000FF0000040404040404040400000000FFFFFFFF0F0F0F0F0F0F0F0F",
		INIT_0F => X"00000000000000FF0101010101010101000000000000FFFF0303030303030303",
		INIT_10 => X"1008080408081000081C3E7F7F1C3E00FF7F3F1F0F070301FFFFFFFFFFFFFFFF",
		INIT_11 => X"081C3663361C0800000010207F2010001C1C6B7F6B081C00003C7E7E7E7E3C00",
		INIT_12 => X"003C424242423C003C42020C10001000FFC381818181C3FF0000000003040808",
		INIT_13 => X"00000000C020101080C0E0F0F8FCFEFF0103070F1F3F7FFF0000080000080000",
		INIT_14 => X"00081C2A080808000E18306030180E003C20202020203C003649414122140800",
		INIT_15 => X"3C04040404043C001C224A564C201E00FFFEFCF8F0E0C08070180C060C187000",
		INIT_16 => X"000808082A1C08000040201008040200000004027F020400F0F0F0F00F0F0F0F",
		INIT_17 => X"000000000F08080800000000F808080808080808F808080800000000FF080808",
		INIT_18 => X"0000013E541414000808080800000800242424000000000024247E247E242400",
		INIT_19 => X"081E281C0A1C08000062640810264600304848304A443A000408100000000000",
		INIT_1A => X"040810101008040020100808081020000008083E08080000082A1C3E1C2A0800",
		INIT_1B => X"0F0F0F0FF0F0F0F08142241818244281101020C0000000000808040300000000",
		INIT_1C => X"FF000000000000008080808080808080FF80808080808080FF01010101010101",
		INIT_1D => X"0000FF0000000000202020202020202001020408102040808040201008040201",
		INIT_1E => X"00000000FF0000000808080808080808FFFFFFFF00000000F0F0F0F0F0F0F0F0",
		INIT_1F => X"000000000000FF0002020202020202020000000000FFFFFF0707070707070707",
		INIT_20 => X"1818181818181800000038043C443A0040405C6242625C0000003C4240423C00",
		INIT_21 => X"02023A4642463A0000003C427E403C000C12107C1010100000003A46463A023C",
		INIT_22 => X"40405C62424242000800180808081C0004000C04040444384040444850684400",
		INIT_23 => X"1808080808081C00000076494949490000005C624242420000003C4242423C00",
		INIT_24 => X"00005C62625C404000003A46463A020200005C624040400000003E403C027C00",
		INIT_25 => X"10107C1010120C000000424242463A0000004242422418000000414949493600",
		INIT_26 => X"000044281028440000004242463A023C00007E0418207E00240038043C443A00",
		INIT_27 => X"0000000102040810031C608000000000C0380601000000000000008040201008",
		INIT_28 => X"00000000C0300C0300FF000000FF0000444444444444444444FF444444FF4444",
		INIT_29 => X"2010080000000000000000324C000000AA44AA11AA44AA1100000000030C30C0",
		INIT_2A => X"030C30C000000000C0300C03000000003844444A42524C000022002222261A00",
		INIT_2B => X"0022001C22221C004200424242423C00421824427E4242004218244242241800",
		INIT_2C => X"1020204040408080010618202040408080601804040202010804040202020101",
		INIT_2D => X"8080404040202010804040202018060101020204041860800101020202040408",
		INIT_2E => X"10080402010000000000000080601C0300000000010638C00810204080000000",
		INIT_2F => X"081010201010080008080808FF08080808142200000000000000000000007E00",
		INIT_30 => X"1C1C3E1C08003E00FFF7F7F7C1E3F7FFFFF7E3C1F7F7F7FFFFFFF7F301F3F7FF",
		INIT_31 => X"FFFFEFCF80CFEFFFBDBDBD81BDBDBDFFE3DDBFBFBFDDE3FF18247EFF5A240000",
		INIT_32 => X"E047427E4247E000223E2A0808497F411C1C083E080814220011D2FCD2110000",
		INIT_33 => X"00884B3F4B880000221408083E081C1C3C7EFFDBFFE77E3C3C4281A58199423C",
		INIT_34 => X"AA55AA55AA55AA550A050A050A050A05A050A050A050A050AA55AA5500000000",
		INIT_35 => X"00000000AA55AA55AA54A850A0408000AA552A150A0502018040A050A854AA55",
		INIT_36 => X"000102050A152A55808040402020101008080404020201013828380000000000",
		INIT_37 => X"00542A542A542A000101020204040808101020204040808000C0C85454552200",
		INIT_38 => X"000000000002FF020202020202020702020202020202FF020000205088050200",
		INIT_39 => X"000E1122C40402011122448811224488007088442320408000C4A4948F94A4C4",
		INIT_3A => X"00232529F12925238890A0C0C0A898B8A8B0B8C0C0A09088804020101F204080",
		INIT_3B => X"00002424E724240008083E00003E0808081020100804020455AA55AA55AA55AA",
		INIT_3C => X"0000000000000000007070700000000000070707000000000077777700000000",
		INIT_3D => X"0000000000707070007070700070707000070707007070700077777700707070",
		INIT_3E => X"0000000000070707007070700007070700070707000707070077777700070707",
		INIT_3F => X"0000000000777777007070700077777700070707007777770077777700777777",
		INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
	port map (
      DOA => D0,      -- Port A 8-bit Data Output
      DOB => CPYD0,      -- Port B 8-bit Data Output
      DOPA => open,    -- Port A 1-bit Parity Output
      DOPB => open,    -- Port B 1-bit Parity Output
      ADDRA => XA,  -- Port A 11-bit Address Input
      ADDRB => CPYA,  -- Port B 11-bit Address Input
      CLKA => DCLK,    -- Port A Clock
      CLKB => PCGDSEL,    -- Port B Clock
      DIA => net_gnd,      -- Port A 8-bit Data Input
      DIB => net_gnd,      -- Port B 8-bit Data Input
      DIPA => net_gnd(0 downto 0),    -- Port A 1-bit parity Input
      DIPB => net_gnd(0 downto 0),    -- Port-B 1-bit parity Input
      ENA => net_vcc,      -- Port A RAM Enable Input
      ENB => net_vcc,      -- PortB RAM Enable Input
      SSRA => net_gnd(0),    -- Port A Synchronous Set/Reset Input
      SSRB => net_gnd(0),    -- Port B Synchronous Set/Reset Input
      WEA => net_gnd(0),      -- Port A Write Enable Input
      WEB => net_gnd(0)       -- Port B Write Enable Input
	);

	--
	-- RAM (CG data included:alternate)
	--
   RAMB16_S9_S9_inst1 : RAMB16_S9_S9
	generic map (
      INIT_A => X"000", --  Value of output RAM registers on Port A at startup
      INIT_B => X"000", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"000", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"000", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "READ_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "READ_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
		INIT_00 => X"00000000000000007C82BABA82BAAAEEFC86BA84BABA86FC7E82BEA0A0BE827E",
		INIT_01 => X"F886B6AAAAB686F8FE82BE8888BE82FEFE82BE88B8A0A0E07E82BEA0AEBA827E",
		INIT_02 => X"EEAABA82BAAAAAEEFE82EE2828EE82FE1F111B0AEABAC67CE6AAB48888B4AAE6",
		INIT_03 => X"E0A0A0A0A0BE82FEFE82AAAABAAAAAEEEE9A8AA2B2AAAAEE7CC6BAAAAABAC67C",
		INIT_04 => X"FC86BABA86BCA0E07CC6BABAAAB2C27CFC86BABA84B4AAE67EC2BEC47AFA86FC",
		INIT_05 => X"FE82EE2828282838EEAAAAAAAABAC67CEEAAAAAAAA542810EEAAAABAAAAA82FE",
		INIT_06 => X"C6AA54282854AAC6EEAA924428282838FE82FA14285E82FE0040A090FF7E0000",
		INIT_07 => X"00020509FF7E0000007CD67C38549200925438FE3854920000003854FE000000",
		INIT_08 => X"7C82B2AAAA9A827C38486828286C447C7C82BACA142E42FEFC82FA2222FA82FC",
		INIT_09 => X"0C142454B682F61CFE82BE847AFA86FC7E82BEBC82BA827CFE82FA1428505070",
		INIT_0A => X"7C82BA7C82BA827C7C82BA827AFA82FCF888BEAAFA223E001F117D555F447C00",
		INIT_0B => X"3C5AFFE77E2442813C5AFFE77E242466081C2A7F773E3663081C2A7F773E3614",
		INIT_0C => X"41A23C5A7EFF426382453C5A7EFF42C6005ABD992442240081A55A181824C300",
		INIT_0D => X"00247EBD7E2424E7247EBD7E244242C33C5AFFABD5FFDD893C5AFFABD5FF7722",
		INIT_0E => X"3C42A5819981D5AA3C42A5819981AB55424266E7FFFF7E3C1CFE3F0F0F3FFE1C",
		INIT_0F => X"3C7EFFFFE7664242387FFCF0F0FC7F383C7EFFFFFFFF7E3C10382828287CFED6",
		INIT_10 => X"0003077EC77E07036B7F3E1414141C0800C0E07EE37EE0C03C0C3C183C767646",
		INIT_11 => X"3C243C183C5A5A7E3C303C183C6E6E627E7E24242424246C7E7E242424242466",
		INIT_12 => X"7E7E2424242424362263F7B7FF7E3C3C386CFF3F0F3FFC383C3C7EFFEDEFC644",
		INIT_13 => X"1C36FFFCF0FC3F1E3C7EFFBFFF7E3C3C3C3C7EFFFDFF7E3C1C36FFFFFFFF3E1C",
		INIT_14 => X"386CFFFFFFFF7C38183C3C3C3C183C3C00007BFFFF7B00003C3C183C3C3C3C18",
		INIT_15 => X"0000DEFFFFDE00002060202030283C3C0040FF0B070300003C3C140C04040604",
		INIT_16 => X"0002FFD0E0C000001010387C9210103800081031FF311008381010927C381010",
		INIT_17 => X"0010088CFF8C081000786050480402000002044850607800004020120A061E00",
		INIT_18 => X"001E060A12204000187E7EFFC38181811F7870F0F070781F818181C3FF7E7E18",
		INIT_19 => X"F81E0E0F0F0E1EF8BFA1ADA5A5BD81FFFF81BDA585FD01FFFF81BDA5A5B585FD",
		INIT_1A => X"FF80BFA1A5BD81FF0018003C007E00FF0105155555150501FF007E003C001800",
		INIT_1B => X"80A0A8AAAAA8A08000081C3E00081C3E0000113377331100003E1C08003E1C08",
		INIT_1C => X"00004466776644000000E7A5E7000000103854101054381000002442FF422400",
		INIT_1D => X"7F41221C0808087F5555555555555555FF00FF00FF00FF00A542A50000A542A5",
		INIT_1E => X"2442810000814224FF809FA0A0A0A0A0FF01E51115111511000000FFA0AFA0FF",
		INIT_1F => X"000000FF414155FFA09F80FF3030307811E101FF0C0C0C1E80AA8095808F80FF",
		INIT_20 => X"01A9015101E101FF3C42ABD51010140800001824241800000018244242241800",
		INIT_21 => X"3C4281818181423C000000181800000000003C3C3C3C0000007E7E7E7E7E7E00",
		INIT_22 => X"3C429DA1A19D423CFFFFFFE7E7FFFFFFFFFFC3C3C3C3FFFFFF818181818181FF",
		INIT_23 => X"20302020FF7E3C003C4281FFFF81423C3C5A999999995A3C3C5A99FFFF995A3C",
		INIT_24 => X"0028FEAAFE5438100F30404E8A8E8081F00C0272517101810F3040408E808081",
		INIT_25 => X"F00C020271010181818088844340300F81011121C2020CF0818080874040300F",
		INIT_26 => X"810101E102020CF0818083844340300F8101C121C2020CF0818087884840300F",
		INIT_27 => X"8101E11112020CF0081054FEFEFEFE7C000608103078783000523406602C4A00",
		INIT_28 => X"91520003C0004A8980C0E0F0FFFFFFFF00000102FFC3C3FF00008040FFC3C3FF",
		INIT_29 => X"00C02010FCFEFFFC0103070FFFFFFFFF021428081414080000FE4220102042FE",
		INIT_2A => X"000304083F7FFF3F0020101010284886003C42424224A5E700448282926C0000",
		INIT_2B => X"00006C92926C000000026C90906E0000001E105050B01000000010007C001000",
		INIT_2C => X"00F15B5555515100FF8991C5A38991FFFFC3A59999A5C3FF00925438EE385492",
		INIT_2D => X"FF9999FFFF9999FF92543810101010103810381038103810000000AAFFAA0000",
		INIT_2E => X"0010107C1010007C7E427E427E427E4200FF55555555FF00000000C0B08C83FF",
		INIT_2F => X"000000030D31C1FF000000003C7EFFFFFFFF7E3C00000000C0E0F0F0F0F0E0C0",
		INIT_30 => X"03070F0F0F0F0703030C3F3FFF7F371FC030B8DCEEF6FBFB0E0E0A040101030F",
		INIT_31 => X"7A74F4F4F4FAFDFD044EE4466F7F603F20722762F6FE06FC3B311B1F101F0F07",
		INIT_32 => X"DC8CD8F808F8F0E0010307060E3E703080C0E060707C0E0C1E0E060703377F8B",
		INIT_33 => X"787060E0C0ECFED101337B598CDF7F3F80CCDE9A31FBFEFC3F1F1F0F0F7F00FF",
		INIT_34 => X"FCF8F8F0F0FE00FF0001020402011F1F008040204080F8F8020202021F207F00",
		INIT_35 => X"40404040F804FE007373737F3F1F0F0FCECECEFEFCF8F0F00F0F0F187F407FFF",
		INIT_36 => X"F0F0F018FE02FEFFF8444221214244F8FF050700000705FFFC868281818286FC",
		INIT_37 => X"000080407F80000000000000FF01010101010101FF000000FF80808080000000",
		INIT_38 => X"00000000808080FF00080C0AF90A0C0800080C3AE93A0C081F2848FE88888F00",
		INIT_39 => X"40C040E60902040F40C040E2060A1F0240C040EF0107010F40A0204FE107010F",
		INIT_3A => X"C0601806186080FE010618601806017F0001061D2A2A2A1F1B8F6511C9A9B1F3",
		INIT_3B => X"4CF7F01807023EFE7F9F31418181F9FD88024000884100914001880040048011",
		INIT_3C => X"003058FDFF793000000C1ABFFF9E0C00003058FD3FF93000000C1ABFFC9F0C00",
		INIT_3D => X"102868BCFC781038BAEEAA3838BAFEBABAFEBA3838AAEEBA00E742FF9FFF42E7",
		INIT_3E => X"00E742FFF9FF42E70000FC1C7F633E0000003F38FEC67C00FF81A58181A581FF",
		INIT_3F => X"E7818100008181E7000408FE10FE204018242420101010100808080804242418",
		INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
	port map (
      DOA => D1,      -- Port A 8-bit Data Output
      DOB => CPYD1,      -- Port B 8-bit Data Output
      DOPA => open,    -- Port A 1-bit Parity Output
      DOPB => open,    -- Port B 1-bit Parity Output
      ADDRA => XA,  -- Port A 11-bit Address Input
      ADDRB => CPYA,  -- Port B 11-bit Address Input
      CLKA => DCLK,    -- Port A Clock
      CLKB => PCGDSEL,    -- Port B Clock
      DIA => net_gnd,      -- Port A 8-bit Data Input
      DIB => net_gnd,      -- Port B 8-bit Data Input
      DIPA => net_gnd(0 downto 0),    -- Port A 1-bit parity Input
      DIPB => net_gnd(0 downto 0),    -- Port-B 1-bit parity Input
      ENA => net_vcc,      -- Port A RAM Enable Input
      ENB => net_vcc,      -- PortB RAM Enable Input
      SSRA => net_gnd(0),    -- Port A Synchronous Set/Reset Input
      SSRB => net_gnd(0),    -- Port B Synchronous Set/Reset Input
      WEA => net_gnd(0),      -- Port A Write Enable Input
      WEB => net_gnd(0)       -- Port B Write Enable Input
	);

	--
	-- RAM (PCG data area)
	--
   RAMB16_S9_S9_inst2 : RAMB16_S9_S9
   generic map (
      INIT_A => X"000", --  Value of output RAM registers on Port A at startup
      INIT_B => X"000", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"000", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"000", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "READ_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "READ_FIRST") --  WRITE_FIRST, READ_FIRST or NO_CHANGE
   port map (
      DOA => D2,      -- Port A 8-bit Data Output
      DOB => open,      -- Port B 8-bit Data Output
      DOPA => open,    -- Port A 1-bit Parity Output
      DOPB => open,    -- Port B 1-bit Parity Output
      ADDRA => EXA,  -- Port A 11-bit Address Input
      ADDRB => PCGA,  -- Port B 11-bit Address Input
      CLKA => DCLK,    -- Port A Clock
      CLKB => PCGWP,    -- Port B Clock
      DIA => net_gnd,      -- Port A 8-bit Data Input
      DIB => PCGD,      -- Port B 8-bit Data Input
      DIPA => net_gnd(0 downto 0),    -- Port A 1-bit parity Input
      DIPB => net_gnd(0 downto 0),    -- Port-B 1-bit parity Input
      ENA => net_vcc,      -- Port A RAM Enable Input
      ENB => net_vcc,      -- PortB RAM Enable Input
      SSRA => net_gnd(0),    -- Port A Synchronous Set/Reset Input
      SSRB => net_gnd(0),    -- Port B Synchronous Set/Reset Input
      WEA => net_gnd(0),      -- Port A Write Enable Input
      WEB => net_vcc       -- Port B Write Enable Input
   );

end Behavioral;
